//write a 4 bit priority counter 
//truth table
//   inputs       output
//  p3 p2 p1 p0   y
//  0  0  0  0    0
//  1  0  0  0    p3
//  0  1  0  0    p2
//  0  0  1  0    p1
//  0  0  0  1    p0

module priority_counter;
  inputs
  outputs

  design code

endmodule
